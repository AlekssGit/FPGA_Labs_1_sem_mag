library verilog;
use verilog.vl_types.all;
entity Lab_4_vlg_vec_tst is
end Lab_4_vlg_vec_tst;
