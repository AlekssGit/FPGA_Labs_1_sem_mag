library verilog;
use verilog.vl_types.all;
entity summ_mod_11_vlg_vec_tst is
end summ_mod_11_vlg_vec_tst;
